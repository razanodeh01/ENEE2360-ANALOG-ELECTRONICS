* C:\Users\Support\NewSemester\Elctro\Project\Part2\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Jul 15 14:03:47 2023



** Analysis setup **
.tran 1m 5m 0 1m
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
